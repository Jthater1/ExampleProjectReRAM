* NGSPICE file created from 1T1R.ext - technology: sky130B

.subckt sky130_fd_pr_reram__reram_cell TE BE
X0 TE BE sky130_fd_pr__reram_reram_cell area_ox=1
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_9YEQ2B a_50_n700# a_n242_n922# a_n108_n700# a_n50_n788#
X0 a_50_n700# a_n50_n788# a_n108_n700# a_n242_n922# sky130_fd_pr__nfet_g5v0d10v5 ad=2.03 pd=14.6 as=2.03 ps=14.6 w=7 l=0.5
.ends

.subckt x1T1R SL VSS WL BL
XXR1 BL XR1/BE sky130_fd_pr_reram__reram_cell
XXM1 XR1/BE VSS SL WL sky130_fd_pr__nfet_g5v0d10v5_9YEQ2B
.ends

