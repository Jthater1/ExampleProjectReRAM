magic
tech sky130B
timestamp 1698708124
<< locali >>
rect 312 -28 340 882
rect 570 -28 598 882
rect 312 -76 598 -28
rect 312 -135 443 -76
rect 591 -135 598 -76
rect 312 -164 598 -135
<< viali >>
rect 443 -135 591 -76
<< metal1 >>
rect 391 462 396 488
rect 425 462 430 488
rect 446 63 466 814
rect 429 36 434 63
rect 479 36 484 63
rect 312 -76 598 -27
rect 312 -135 443 -76
rect 591 -135 598 -76
rect 312 -164 598 -135
<< via1 >>
rect 396 462 425 488
rect 434 36 479 63
<< metal2 >>
rect 347 865 447 965
rect 476 865 576 965
rect 383 488 428 865
rect 383 462 396 488
rect 425 462 428 488
rect 383 461 428 462
rect 396 457 425 461
rect 490 443 535 865
rect 256 56 356 120
rect 434 63 479 68
rect 256 36 434 56
rect 256 32 479 36
rect 256 20 356 32
rect 434 31 479 32
use sky130_fd_pr__nfet_g5v0d10v5_9YEQ2B  XM1
timestamp 1698708124
transform 1 0 455 0 1 427
box -139 -479 139 479
use sky130_fd_pr_reram__reram_cell  XR1
timestamp 1698708124
transform 1 0 484 0 1 572
box -3 -203 103 -97
<< labels >>
flabel metal1 326 -154 426 -54 0 FreeSans 128 0 0 0 VSS
port 1 nsew
flabel metal2 256 20 356 120 0 FreeSans 128 0 0 0 WL
port 2 nsew
flabel metal2 347 865 447 965 0 FreeSans 128 0 0 0 SL
port 0 nsew
flabel metal2 476 865 576 965 0 FreeSans 128 0 0 0 BL
port 3 nsew
<< end >>
